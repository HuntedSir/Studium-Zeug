`timescale 1ns / 1ns

/* ====================================== INSERT CODE HERE ====================================== */

module xor #(SIZE = 2) (
    input logic [SIZE - 1: 0] I,
    output logic O
);

assign O = ^I;
    
endmodule

/* ============================================================================================== */
