`timescale 1ns / 1ns

module comparison #(parameter N)
                  ( input  logic [N-1:0] A, B,
                    output logic         Y);

/* ====================================== INSERT CODE HERE ====================================== */



/* ============================================================================================== */

endmodule

