`timescale 1 ns / 10 ps

module timing_tb;

  //********************* MODULE INPUTS ***********************//
  logic        CLK, R, X, Y;
  //***********************************************************//


  //********************* MODULE OUTPUTS **********************//
  logic        A, B, C, D, E, F, G, H;
  logic [15:0] I, J;
  //***********************************************************//

  //******************* UUT INSTANTIATION *********************//
  timing  uut (CLK, R, X, Y, A, B, C, D, E, F, G, H, I, J);
  //***********************************************************//

  //********************** CLOCK SIGNAL ***********************//
  always begin
    #5 CLK = ~CLK;
  end
  //***********************************************************//

  //********************* TEST INITIATION *********************//
  initial begin
    $dumpfile("timing_tb.vcd");
    $timeformat(-9, 0, " ns", 8);
    $dumpvars;

    CLK = 0;
    X = 1;
    Y = 1;
    R = 1;
    #3;
    X = 0;
    R = 0;
    #4;
    X = 1;
    #1;
    Y = 0;
    #5;
    X = 0;
    #2;
    Y = 1;
    #2;
    X = 1;
    #6;
    Y = 0;
    #4;
    X = 0;
    #1;
    Y = 1;
    #4;
    Y = 0;
    #5;
    X = 1;
    #5;
    Y = 1;
    #1;
    X = 0;
    #4;
    X = 1;
    #5;
    Y = 0;
    #1;
    X = 0;
    #6;
    X = 1;
    #1;
    X = 0;
    #2;
    X = 1;
    Y = 1;
    #1;
    X = 0;
    Y = 0;
    #1;
    X = 1;
    Y = 1;
    #1;
    Y = 0;
    #2;
    Y = 1;
    #6;
    X = 0;
    #1;
    Y = 0;
    #3;
    Y = 1;
    #1;
    X = 1;
    #3;
    Y = 0;
    #2;
    X = 0;
    #1;
    Y = 1;
    #3;
    X = 1;
    #3;
    X = 0;
    #1;
    Y = 0;
    #2;
    X = 1;
    #5;
    Y = 1;
    #2;
        
    $finish;
  end

  //***********************************************************//

endmodule
